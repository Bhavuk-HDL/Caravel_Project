VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO seven_segment_seconds
  CLASS BLOCK ;
  FOREIGN seven_segment_seconds ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 225.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 86.000 55.800 90.000 56.400 ;
    END
  END clk
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 221.000 6.350 225.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 221.000 16.010 225.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 221.000 25.670 225.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 221.000 35.330 225.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 221.000 44.990 225.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 221.000 54.650 225.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 221.000 64.310 225.000 ;
    END
  END io_oeb[6]
  PIN led_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 221.000 73.970 225.000 ;
    END
  END led_out[0]
  PIN led_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END led_out[1]
  PIN led_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END led_out[2]
  PIN led_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END led_out[3]
  PIN led_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 221.000 83.630 225.000 ;
    END
  END led_out[4]
  PIN led_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 86.000 168.000 90.000 168.600 ;
    END
  END led_out[5]
  PIN led_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 4.000 ;
    END
  END led_out[6]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.590 10.640 16.190 212.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.330 10.640 35.930 212.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.070 10.640 55.670 212.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.810 10.640 75.410 212.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.460 10.640 26.060 212.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.200 10.640 45.800 212.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.940 10.640 65.540 212.400 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 84.180 212.245 ;
      LAYER met1 ;
        RECT 5.520 10.640 87.790 212.400 ;
      LAYER met2 ;
        RECT 6.630 220.720 15.450 221.000 ;
        RECT 16.290 220.720 25.110 221.000 ;
        RECT 25.950 220.720 34.770 221.000 ;
        RECT 35.610 220.720 44.430 221.000 ;
        RECT 45.270 220.720 54.090 221.000 ;
        RECT 54.930 220.720 63.750 221.000 ;
        RECT 64.590 220.720 73.410 221.000 ;
        RECT 74.250 220.720 83.070 221.000 ;
        RECT 83.910 220.720 87.760 221.000 ;
        RECT 6.080 4.280 87.760 220.720 ;
        RECT 6.080 4.000 10.850 4.280 ;
        RECT 11.690 4.000 33.390 4.280 ;
        RECT 34.230 4.000 55.930 4.280 ;
        RECT 56.770 4.000 78.470 4.280 ;
        RECT 79.310 4.000 87.760 4.280 ;
      LAYER met3 ;
        RECT 4.000 169.000 86.875 212.325 ;
        RECT 4.000 167.600 85.600 169.000 ;
        RECT 4.000 113.240 86.875 167.600 ;
        RECT 4.400 111.840 86.875 113.240 ;
        RECT 4.000 56.800 86.875 111.840 ;
        RECT 4.000 55.400 85.600 56.800 ;
        RECT 4.000 10.715 86.875 55.400 ;
      LAYER met4 ;
        RECT 31.575 12.415 33.930 111.345 ;
        RECT 36.330 12.415 43.800 111.345 ;
        RECT 46.200 12.415 53.670 111.345 ;
        RECT 56.070 12.415 63.540 111.345 ;
        RECT 65.940 12.415 73.410 111.345 ;
        RECT 75.810 12.415 77.905 111.345 ;
  END
END seven_segment_seconds
END LIBRARY

