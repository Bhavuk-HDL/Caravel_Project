VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO seven_segment_seconds
  CLASS BLOCK ;
  FOREIGN seven_segment_seconds ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 250.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END clk
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 246.000 5.890 250.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 246.000 16.930 250.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 246.000 27.970 250.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 246.000 39.010 250.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 246.000 50.050 250.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 246.000 61.090 250.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 246.000 72.130 250.000 ;
    END
  END io_oeb[6]
  PIN led_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END led_out[0]
  PIN led_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 246.000 83.170 250.000 ;
    END
  END led_out[1]
  PIN led_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END led_out[2]
  PIN led_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 124.480 100.000 125.080 ;
    END
  END led_out[3]
  PIN led_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END led_out[4]
  PIN led_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 246.000 94.210 250.000 ;
    END
  END led_out[5]
  PIN led_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END led_out[6]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.840 10.640 17.440 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.080 10.640 39.680 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.320 10.640 61.920 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.560 10.640 84.160 236.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 26.960 10.640 28.560 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.200 10.640 50.800 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.440 10.640 73.040 236.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 94.300 236.725 ;
      LAYER met1 ;
        RECT 5.520 10.640 94.300 236.880 ;
      LAYER met2 ;
        RECT 6.170 245.720 16.370 246.570 ;
        RECT 17.210 245.720 27.410 246.570 ;
        RECT 28.250 245.720 38.450 246.570 ;
        RECT 39.290 245.720 49.490 246.570 ;
        RECT 50.330 245.720 60.530 246.570 ;
        RECT 61.370 245.720 71.570 246.570 ;
        RECT 72.410 245.720 82.610 246.570 ;
        RECT 83.450 245.720 93.650 246.570 ;
        RECT 5.620 4.280 94.200 245.720 ;
        RECT 5.620 3.670 16.370 4.280 ;
        RECT 17.210 3.670 49.490 4.280 ;
        RECT 50.330 3.670 82.610 4.280 ;
        RECT 83.450 3.670 94.200 4.280 ;
      LAYER met3 ;
        RECT 4.000 208.440 96.000 236.805 ;
        RECT 4.400 207.040 96.000 208.440 ;
        RECT 4.000 125.480 96.000 207.040 ;
        RECT 4.400 124.080 95.600 125.480 ;
        RECT 4.000 42.520 96.000 124.080 ;
        RECT 4.400 41.120 96.000 42.520 ;
        RECT 4.000 10.715 96.000 41.120 ;
      LAYER met4 ;
        RECT 17.840 85.855 26.560 148.745 ;
        RECT 28.960 85.855 37.680 148.745 ;
        RECT 40.080 85.855 48.800 148.745 ;
        RECT 51.200 85.855 59.920 148.745 ;
        RECT 62.320 85.855 71.040 148.745 ;
        RECT 73.440 85.855 76.065 148.745 ;
  END
END seven_segment_seconds
END LIBRARY

